`default_nettype none

module EPP(
    input clk
);


endmodule